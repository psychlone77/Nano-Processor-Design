library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity HA is
    Port ( A : in STD_LOGIC;
           B : in STD_LOGIC;
           C : out STD_LOGIC;
           S : out STD_LOGIC);
end HA;

architecture Behavioral of HA is

begin

C <= A AND B;
--S <= (NOT(A) AND B) OR ((NOT B) AND A);
S <= A XOR B;

end Behavioral;